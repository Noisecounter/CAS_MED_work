-----------------------------------------------------
-- Project : system
-----------------------------------------------------
-- File    : system_top_pkg.vhd
-- Library : system_tb_lib
-- Author  : michael.pichler@fhnw.ch
-- Company : FHNW - ISE
-- Copyright(C) ISE
-----------------------------------------------------
-- Description :
-----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;
use ieee.std_logic_textio.all;

package system_top_pkg is
    -- -------------------------------------------------------
    -- Global Constants & Types
    -- -------------------------------------------------------
    constant C_DWIDTH   : integer := 8;
    constant C_AWIDTH   : natural := 10;
    -- -------------------------------------------------------
    -- Procedure to read data from a memory
    -- -------------------------------------------------------

end system_top_pkg;

package body system_top_pkg is
    -- -------------------------------------------------------
    -- Procedure to read data from a memory
    -- -------------------------------------------------------

end system_top_pkg;
