LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE constants IS
CONSTANT c_max1_syn: integer := 124999;
CONSTANT c_max2_syn: integer := 9;

CONSTANT c_max1_sim: integer := 4;
CONSTANT c_max2_sim: integer := 4;

END constants;


PACKAGE BODY constants IS

END constants;